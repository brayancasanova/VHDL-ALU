library verilog;
use verilog.vl_types.all;
entity test_ALU_vlg_vec_tst is
end test_ALU_vlg_vec_tst;
